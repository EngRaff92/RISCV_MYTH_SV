
module rv32i_core (
	input clk,    			// Clock
	input clk_en, 			// Clock Enable
	input rst,    			// Asynchronous reset active high
`ifdef RV32I_DEBUG	
	output [31:0] pc_debug	// debug Program Counter
`endif
);

	/** Internal signals */
	logic 			gated_clock;
    logic [31:0]  	core_in_branch;
    logic [31:0]  	core_in_jump;
    logic         	core_is_jump;
    logic         	core_is_branch;
`ifdef RV32I_DEBUG	    
    logic [31:0] 	core_pc;
    logic           core_r_type_instr_o;
    logic           core_i_type_instr_o;
    logic           core_s_type_instr_o;
    logic           core_b_type_instr_o;
    logic           core_u_type_instr_o;
    logic           core_j_type_instr_o;
    logic           core_illegal_instr_o;
    logic [2:0]     core_funct3_o;
`endif    
    logic        	core_pc_error;
    logic [31:0]	core_instr_i;
    logic [4:0]     core_rs1_o;
    logic [4:0]     core_rs2_o;
    logic [4:0]     core_rd_o;
    logic [6:0]     core_op_o;
    logic [6:0]     core_alu_op_sel_0;
    logic [19:0]    core_instr_imm_;
  	logic [31:0]    core_opr_a_i;		
  	logic [31:0]    core_opr_b_i;
  	logic [31:0] 	core_alu_res_o;
	logic [3:0]  	core_op_sel_i;
	logic 			core_rf_cs;
	logic 			core_d_cs;
	logic [9:0] 	core_mem_addr;
	
	/** Gating cell */
	clock_g u_clock_gating_cell(
		.clk_en   (clk_en),	
		.clk_in   (clk),
		.clock_out(gated_clock));

	/** Instruction Uunit */
	instruction_fetch u_fecth_unit(
		.fetch_rst 			(rst),
		.fetch_clk 			(gated_clock),
		.in_branch 			(core_in_branch),
		.in_jump  			(core_in_jump),
		.is_jump  			(core_is_jump),
		.is_branch 			(core_is_branch),
`ifdef RV32I_DEBUG
		.pc       			(core_pc),
`endif
		.instruction_fecthed(core_instr_i),
		.pc_error 			(core_pc_error));

	/** Decoder Unit */
	opcode_decoder u_decoder_unit(
		.instr_i        (core_instr_i),
		.rs1_o          (core_rs1_o),
		.rs2_o          (core_rs2_o),
		.rd_o           (core_rd_o),
		.op_o           (core_op_o),			
		.alu_op_sel_0   (core_alu_op_sel_0),	/** ALU operation using func7 + func5*/
`ifdef RV32I_DEBUG		
		.funct3_o       (core_funct3_o),		/** func3 used by the control unit to detect the Instruction type */
		.r_type_d 		(core_r_type_instr_o),
		.i_type_d 		(core_i_type_instr_o),
		.s_type_d 		(core_s_type_instr_o),
		.b_type_d 		(core_b_type_instr_o),
		.u_type_d 		(core_u_type_instr_o),
		.j_type_d 		(core_j_type_instr_o),
		.illegal_d 		(core_illegal_instr_o),
`endif
		.instr_imm_o    (core_instr_imm_o),  	/** immediate generated by the immedaite unit */
		.memory_address (core_mem_addr));

	/** Control Unit */
	opcode_control_unit u_control_unit(
		.in_intruction  (in_intruction),
		.reg_file_w_r_en(reg_file_w_r_en),
		.memory_r_w_en  (memory_r_w_en),
		.reg_file_cs    (reg_file_cs),
		.memory_cs      (memory_cs),
		.write_back     (write_back),
		.memory_address (memory_address));

	/** Register file Unit */
	register_file u_register_file(
		.rf_clk   (gated_clock),
		.rf_ares  (rst),
		.rw_dec   (core_rd_o),
		.ra_dec   (core_rs1_o),
		.rb_dec   (core_rs2_o),
		.w_data_in(core_alu_res_o),
		.rf_cs	  (core_rf_cs),
		.wr_en    (core_r_type_instr_o),
		.qa_out   (core_opr_a_i),
		.qb_out   (core_opr_b_i));

	/** Alu Unit */
	rv_alu u_alu_unit(
		.opr_a_i  (core_opr_a_i),
		.opr_b_i  (core_opr_b_i),
		.op_sel_i (core_alu_op_sel_0),
		.alu_res_o(core_alu_res_o));

	/** Data memory Unit */
	data_memory#(10,10,32,0) u_data_memory_unit(
		.d_clk   (clk),
		.d_rst   (rst),
		.d_addr  (core_mem_addr),
		.d_w_data(d_w_data),
		.d_cs    (core_d_cs),
		.d_rw_en (d_rw_en),
		.d_r_data(d_r_data));

`ifdef RV32I_DEBUG
	/** Assign the debug programm counter */
	assign pc_debug = core_pc;
`endif
endmodule // rv32i_core