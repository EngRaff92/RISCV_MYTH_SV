/** Main Write Back unit */

module write_back_unit(
	// Input ports
	input logic write_back_enable);

	/** Main */
endmodule // write_back_unit