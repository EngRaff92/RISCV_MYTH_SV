
module rv32i_core (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
);

endmodule // rv32i_core